module lcd_driver(
	
);
